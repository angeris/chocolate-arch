module regfile(
    
)